LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SELECIONA_DESTINO IS
	port(
		i_CLK 					: IN STD_LOGIC;
		i_RST						: IN STD_LOGIC;
		i_DESTINO_E				: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		i_DESTINO_D				: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		i_CONFIRMA_E			: IN STD_LOGIC;
		i_CONFIRMA_D			: IN STD_LOGIC;
		i_CONFIRMA_PAINEL_E 	: IN STD_LOGIC;
		i_CONFIRMA_PAINEL_D 	: IN STD_LOGIC;
		i_ANDAR_VIAGEM			: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		o_CONFIRMA_E			: OUT STD_LOGIC;
		o_CONFIRMA_D			: OUT STD_LOGIC;
		o_DESTINO_E				: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		o_DESTINO_D				: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);	
END SELECIONA_DESTINO;


ARCHITECTURE BEHAVORIAL OF SELECIONA_DESTINO IS	
BEGIN

	PROCESS(i_CLK, i_RST)
	BEGIN
		if(i_RST = '0') THEN
			o_CONFIRMA_D 	<= '0';
			o_CONFIRMA_E	<= '0';
			o_DESTINO_D 	<= "00";
			o_DESTINO_E		<= "00";
		elsif RISING_EDGE(i_CLK) THEN
			if(i_CONFIRMA_PAINEL_E = '0') THEN
				o_CONFIRMA_E <= i_CONFIRMA_PAINEL_E;
				o_DESTINO_E <= i_ANDAR_VIAGEM;
			else
				o_CONFIRMA_E <= i_CONFIRMA_E;
				o_DESTINO_E <= i_DESTINO_E;
			end if;
			
			if(i_CONFIRMA_PAINEL_D = '0') THEN
				o_CONFIRMA_D <= i_CONFIRMA_PAINEL_D;
				o_DESTINO_D  <= i_ANDAR_VIAGEM;
			else
				o_CONFIRMA_D <= i_CONFIRMA_D;
				o_DESTINO_D <= i_DESTINO_D;
			END IF;
		END IF;
	END PROCESS;
END;


	
	