	LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_ARITH.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_ELEVADOR IS
END TB_ELEVADOR;

ARCHITECTURE BEHAVIORAL OF TB_ELEVADOR IS

	COMPONENT ELEVADOR IS
		port(
					i_CLK								: IN STD_LOGIC;					
					i_RST								: IN STD_LOGIC;
					i_DESTINO						: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
					i_CONFIRMA_NOVO_DESTINO		: IN STD_LOGIC;
					o_PORTAS							: OUT STD_LOGIC;
					o_MOVIMENTO						: OUT STD_LOGIC;
					o_ANDAR_ATUAL					: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
		);
	end COMPONENT;

SIGNAL w_CLK, w_RST, w_CONFIRMA_NOVO_DESTINO : STD_LOGIC;
SIGNAL w_PORTAS, w_MOVIMENTO : STD_LOGIC;
SIGNAL w_ANDAR_ATUAL : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL w_DESTINO : STD_LOGIC_VECTOR(1 DOWNTO 0);

	PROCEDURE CLK_GEN(signal w_CLK : OUT STD_LOGIC; constant FREQ: INTEGER) IS
		CONSTANT PERIOD : time := 1 sec / FREQ;
		BEGIN
			LOOP
				w_CLK <= '1';
				wait for PERIOD/2;
				w_CLK <= '0';
				wait for PERIOD/2;
			END LOOP;
	END PROCEDURE;

BEGIN
	U001 : ELEVADOR
		PORT MAP(
			i_CLK								=> w_CLK,
			i_RST								=> w_RST,
			i_DESTINO						=> w_DESTINO,
			i_CONFIRMA_NOVO_DESTINO		=> w_CONFIRMA_NOVO_DESTINO,
			o_PORTAS							=> w_PORTAS,
			o_MOVIMENTO						=> w_MOVIMENTO,
			o_ANDAR_ATUAL					=> w_ANDAR_ATUAL
		);
	
CLK_GEN(w_CLK, 50000000);

PROCESS
	BEGIN
		w_RST <= '0';
		wait for 200 ns;
		w_RST <= '1';
		wait for 200 ns;
		
		w_DESTINO <= "10";
		w_CONFIRMA_NOVO_DESTINO <= '0';
		
		wait for 5 us;
		
		w_DESTINO <= "00";
		w_CONFIRMA_NOVO_DESTINO <= '0';
		
		wait for 5 us;
	END PROCESS;
END;
		