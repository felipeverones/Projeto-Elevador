	LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_ARITH.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;

	ENTITY TIMER IS
	
	PORT(
		i_CLK				: IN STD_LOGIC;
		i_RST				: IN STD_LOGIC;
		i_EN				: IN STD_LOGIC;
		i_DATA			: IN STD_LOGIC_VECTOR(27 DOWNTO 0); -- 1011 1110 1011 1100 0010 0000 0000 = 4s
		i_RELOAD			: IN STD_LOGIC;
		o_EST				: OUT STD_LOGIC
	);
END TIMER;

ARCHITECTURE BEHAVIORAL OF TIMER IS

SIGNAL w_COUNT : STD_LOGIC_VECTOR(27 DOWNTO 0);

BEGIN

PROCESS(i_CLK, i_RST, i_RELOAD)
	BEGIN
	if(i_RST = '0') THEN
		o_EST <= '0';
	elsif(i_RELOAD = '1') THEN
			w_COUNT <= i_DATA;
			o_EST <= '0';
	elsif RISING_EDGE(i_CLK) THEN
		if(i_EN = '1') THEN
			if(w_COUNT /= "0000000000000000000000000000")THEN
				w_COUNT <= w_COUNT - 1;
				o_EST <= '0';
			elsif(w_COUNT = "0000000000000000000000000000") THEN
				o_EST <= '1';
			end if;
		end if;
	else
	end if;
	END PROCESS;
END;
		